parameter renderH = 240;
parameter renderV = 180;
parameter outputH = 960;
parameter outputV = 640;

parameter hsync = 96;
parameter hbackporch = 136;
parameter hfrontporch = 40;

parameter vsync = 10;
parameter vbackporch = 12;
parameter vfrontporch = 3;

parameter pixelClk = 49; //49 MHz may end up not using