//try to make this pur
module pixel_decoder #(DATA_WIDTH=16) (
    input 
)

endmodule